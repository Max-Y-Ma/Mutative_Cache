interface gpio_itf #(parameter NUM_GPIO = 8);

wire [NUM_GPIO-1:0] gpio;

endinterface
