module mutative_fsm (
    input   logic           clk,
    input   logic           rst,


);


endmodule