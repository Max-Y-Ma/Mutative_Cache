interface adp_itf;

logic       tck;
logic       tms;
logic       tdi;
logic       tdo;
logic [3:0] tst;

endinterface
