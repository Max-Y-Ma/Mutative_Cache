interface uart_itf;

logic tx;
logic rx;

endinterface