interface spi_itf;

logic mosi;
logic miso;
logic cs;
logic sclk;

endinterface
