interface spi_itf;

logic mosi;
logic sclk;

endinterface
