// Configuration for UVM Testbench for RISCV Pipeline CPU
`define NUM_TEST (1000000)
`define NOP_INSTR (32'h13)