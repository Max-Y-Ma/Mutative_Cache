interface i2c_itf;

wire  sda;
logic scl;

endinterface
